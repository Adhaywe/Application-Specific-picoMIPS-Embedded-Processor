//File name: opcodes.sv
//Function: pMIPS opcode definitions

`define NOP 6'b000000
`define IO1 6'b000110
`define IO2 6'b001110
`define ADD 6'b000010
`define ADDI 6'b001010
`define LDI 6'b011010
`define MULTI 6'b000011
`define J 6'b000101





