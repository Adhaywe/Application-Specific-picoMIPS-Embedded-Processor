//File name: alucodes.sv
//Function: pMIPS ALU function code definitions


`define RADD 3'b010
`define RSUB 3'b111
`define RMUL 3'b011
 
